    Mac OS X            	   2  �     �                                    ATTR      �   �   �                  �   �  "com.apple.LaunchServices.OpenWith      a     com.apple.lastuseddate#PS idebplist00�WversionTpath_bundleidentifier _!/System/Applications/TextEdit.app_com.apple.TextEdit/1U                            j�$�g    k�+$                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��