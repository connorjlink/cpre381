-------------------------------------------------------------------------
-- Author: Connor Link
-- Date: 02.11.2025
-- Files: RISCV_types.vhd
-------------------------------------------------------------------------
-- Description: This file contains some types that 3810 students
-- may want to use for their RISC-V implementation. This file is guaranteed to 
-- compile first, so if any types, constants, functions, etc., etc., are wanted, 
-- students should declare them here.
-------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;

package RISCV_types is

-- Generic placeholders to define the bit widths for our architecture
constant DATA_WIDTH : natural := 32;
constant ADDR_WIDTH : natural := 10;

-- Type declaration for the register file storage
type array_t is array (natural range <>) of std_logic_vector(31 downto 0);

-- Corresponding func3 values for each branch type
constant BEQ  : natural := 1;
constant BNE  : natural := 2;
constant BLT  : natural := 3;
constant BGE  : natural := 4;
constant BLTU : natural := 5;
constant BGEU : natural := 6;
constant J    : natural := 7; -- force jump for `jal` and `jalr`

-- Corresponding to each load/store data width
constant BYTE   : natural := 0;
constant HALF   : natural := 1;
constant WORD   : natural := 2;
constant DOUBLE : natural := 3;

-- Corresponding to each ALU operation code input signal
constant ADD  : natural := 0;
constant SUB  : natural := 1;
constant BAND : natural := 2;
constant BOR  : natural := 3;
constant BXOR : natural := 4;
constant BSLL : natural := 5;
constant BSRL : natural := 6;
constant BSRA : natural := 7;
constant SLT  : natural := 8;
constant SLTU : natural := 9;

-- Corresponding to each RF source command
constant FROM_RAM    : natural := 1;
constant FROM_ALU    : natural := 2;
constant FROM_NEXTIP : natural := 3;
constant FROM_IMM    : natural := 4;

-- Corresponding to each branch mode type (for correct effective address calculation)
constant JAL_OR_BCC : natural := 1;
constant JALR       : natural := 2;


-- Record type declarations for the pipeline setup
-- Instruction register -> Driver
type insn_record_t is record
    IPAddr   : std_logic_vector(31 downto 0);
    LinkAddr : std_logic_vector(31 downto 0);
    Insn     : std_logic_vector(31 downto 0);
end record insn_record_t;

-- Driver -> ALU
type driver_record_t is record
    MemWrite   : std_logic;
    RegWrite   : std_logic;
    RFSrc      : natural;
    ALUSrc     : std_logic;
    ALUOp      : natural;
    BGUOp      : natural;
    LSWidth    : natural;
    RD         : std_logic_vector(4 downto 0);
    RS1        : std_logic_vector(4 downto 0);
    RS2        : std_logic_vector(4 downto 0);
    DS1        : std_logic_vector(31 downto 0);
    DS2        : std_logic_vector(31 downto 0);
    Imm        : std_logic_vector(31 downto 0);
    BranchMode : natural;
    nInc2_Inc4 : std_logic;
    IPToALU    : std_logic;
end record driver_record_t;

-- ALU -> Memory
type alu_record_t is record
    F  : std_logic_vector(31 downto 0);
    Co : std_logic;
end record alu_record_t;

-- Memory -> Register file
type mem_record_t is record
    Data : std_logic_vector(31 downto 0);
end record mem_record_t;


end package RISCV_types;

-- package body RISCV_types is
--     -- This section is intentionally left blank
-- end package body RISCV_types;
