    Mac OS X            	   2  �     �                                    ATTR      �   �   �                  �   �  "com.apple.LaunchServices.OpenWith      f     com.apple.lastuseddate#PS idebplist00�WversionTpath_bundleidentifier _$/Applications/Visual Studio Code.app_com.microsoft.VSCode/1X                            o���g    )��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             This resource fork intentionally left blank                                                                                                                                                                                                                            ��